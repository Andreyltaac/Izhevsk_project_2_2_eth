module only_rx (


	input														clk_l, 
	input														clk_h,
	input														clk_hh,
	input														rst,

	input 			[3:0]										ss_in,
	input 			[2:0]										m_in,
	input           [2:0]                                       bw_in,
	input			[23:0]										thr_lvl,
	input			[1:0]										frsync_ctrl,

	input			[15:0]										rx_i_axis_tdata,
	input														rx_i_axis_tvalid,
	output														rx_i_axis_tready,
	input			[15:0]										rx_q_axis_tdata,
	input														rx_q_axis_tvalid,
	output														rx_q_axis_tready,
	input 			[13:0]										addr_shft,
	output     													corr_pr_detect,
	output                                                      DeFec_err_dtct,
	output                                                      decrc_oerr,
	output                                                      decrc_verr,
	output                                                      finder_osop,
	output                                                      p1_verr,
	output                                                      p2_oerr,
	output                                                      time_er,
	output                                                      rx_ocorr_dtct,
	output			[23:0]										delta_ph,
	output          [17:0]                                      kb_ps,
	output			[31:0]			                            corr_sig,


	output			[23:0]										thr_lvl_auto,
	output			[14:0]										N_sop_detect,
	output			[23:0]										N_err,
	output			[7:0]										m_axis_tdata,
	output														m_axis_tvalid,
	output														m_axis_tlast,
	output			[0:0]										m_axis_tuser,
	input														m_axis_tready,

	input														m_axis_aclk,
	input														rx_i_axis_aclk,
	input														rx_q_axis_aclk
);

wire signed [4:0]		phy_fifo_dat;
wire 					phy_fifo_val;
wire signed [7:0]		fifo_defec_dat;
wire 					fifo_defec_val;


assign rx_i_axis_tready = 1'd1;
assign rx_q_axis_tready = 1'd1;

RX_phy
RX_phy_sub(
		.clk_low_data		(clk_l),
		.clk_h				(clk_h),
		.rst				(rst),
		.ss_in				(ss_in),
		.m_in				(m_in),
	    .fr_sync_ctrl		(frsync_ctrl),
		.bw_in				(bw_in),
		.thr_lvl			(thr_lvl),
		.addr_shft			(addr_shft),
		.n_sps				(N_sop_detect),
		.m_ax_obit_soft		(phy_fifo_dat),
		.m_ax_oval_soft		(phy_fifo_val),
		.thr_lvl_auto		(thr_lvl_auto),
		.corr_sig           (corr_sig),
		.corr_pr_detect		(corr_pr_detect),
		.ocorr_dtct         (rx_ocorr_dtct),
		.isub_i				(rx_i_axis_tdata),
		.isub_q				(rx_q_axis_tdata),
		.delta_ph			(delta_ph));


axis_data_fifo_fhy_defec axis_data_fifo_fhy_defec_sub (
  .s_axis_aresetn	(rst), 
  .s_axis_aclk		(clk_h),       
  .s_axis_tvalid	(phy_fifo_val),   
  .s_axis_tready	(),   
  .s_axis_tdata		({3'd0, phy_fifo_dat}),     

  .m_axis_aclk		(clk_hh),       
  .m_axis_tvalid	(fifo_defec_val),   
  .m_axis_tready	(1'd1),   
  .m_axis_tdata		(fifo_defec_dat)      
);

wire	[7:0]		m_axis_tdata_l;
wire				m_axis_tvalid_l;
//wire				decrc_oerr;
 DeFEC DeFEC_sub(
    	.clk			(clk_hh),
    	.rst			(rst),
    	.idat			(fifo_defec_dat[4:0]),
		.ival			(fifo_defec_val),
		.ordy			(),
    	.irdy			(),
    	.oval			(m_axis_tvalid_l),
    	.odat			(m_axis_tdata_l),
		.err_dtct       (DeFec_err_dtct),
		.decrc_verr     (decrc_verr),
		.decrc_oerr		(decrc_oerr),
		.finder_osop    (finder_osop));





wire	odgood, oval_prbs;

prbs23_check
#(
  .pDAT_W			( 8),
  .pMSB_FIRST		( 0),  // 1/0 :: first scrambled bit is MSB/LSB
  .pERR_PERIOD_W	(24),
  .pERR_W			(15))
prbs23_check_sub 
(
  .iclk			(clk_hh),
  .iclkena		(1'd1),
  .ibyp			(1'd0),
  .iclr			(~rst),
  .ival			(m_axis_tvalid_l),
  .idat			(m_axis_tdata_l),
  .oval			(oval_prbs),
  .odat			(),
  .err			(),
  .err_led		(),
  .odgood		(odgood)
);


count_err
count_err_sub(
	.clk	(clk_hh),
	.rst	(~rst),
	.err	(odgood),
	.val	(oval_prbs),
	.n_er	(N_err)
);


assign m_axis_tdata	 =	m_axis_tdata_l;
assign m_axis_tvalid =	m_axis_tvalid_l;
assign m_axis_tlast  =	0;
assign m_axis_tuser	 =  0;


speed_test #(
    .B1(1920)  // �?зменение на 5 единиц
) speed_test_sub 
(
    .clk      (clk_l),
    .clk_hh   (clk_hh),
    .reset    (~rst),
    .p1       (decrc_verr),
    .p2       (decrc_oerr),
    .d1_out   (kb_ps),
    .valid_out(time_er),
	.p1_rise  (p1_verr),
	.p2_rise  (p2_oerr)
);


endmodule